package frame_en_lib;
    `define hsl_v3                      1
endpackage
